`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Create Date: 07/16/2023 01:13:34 PM
// 
//////////////////////////////////////////////////////////////////////////////////

`define reset_all() \
    // Address Write Channel \
    axi_awaddr = 5'b0000; \
    axi_awvalid = 1'b0; \
    // Write Channel \
    axi_wdata = 32'h0000; \
    axi_wstrb = 4'b0000; \
    axi_wvalid = 1'b0; \
    // Write Response Channel \
    axi_bready = 1'b0; \
    // Read Address Channel \
    axi_araddr = 5'b00000; \
    axi_arprot = 3'b000; \
    axi_arvalid = 1'b0; \
    // Read Data Channel \
    axi_rready = 1'b0;

module test_bench(

    );
    
    // Clock Signal 100MHz
    reg clk;
    initial begin
        clk = 0;
        forever #(5) clk = !clk;  //100MHz clock
    end

    wire scl_io; // Read only - slave never drives

    wire sda_io; // Connect to sda_io
    reg sda_drive;
    reg sda_tx;
    assign sda_io = (sda_drive)? sda_tx: 1'bZ;

    wire req_data_chunk;
    wire busy;
    wire nack;

    reg axi_aresetn;

    reg  [ 4:0]  axi_awaddr;
    reg  [ 2:0]  axi_awprot;
    reg          axi_awvalid;
    wire         axi_awready; // output
    
    reg  [31:0]  axi_wdata; 
    reg  [ 3:0]  axi_wstrb;
    reg          axi_wvalid;
    wire         axi_wready; // output

    wire [ 1:0]  axi_bresp; // output
    wire         axi_bvalid; // output
    reg          axi_bready;

    reg  [ 4:0]  axi_araddr;
    reg  [ 2:0]  axi_arprot;
    reg          axi_arvalid;
    wire         axi_arready; // output

    wire [31:0]  axi_rdata; // output
    wire [ 1:0]  axi_rresp; // output
    wire         axi_rvalid; // output
    reg          axi_rready;

    // Local variable for reading results from the I2C/SDA
    reg [7:0] tmp_result;

    // Run Tests Here
    initial begin
        $timeformat(-9, 2, " ns", 20);

        axi_aresetn = 0;
        sda_drive = 0;
        `reset_all

        #50;
        axi_aresetn = 1;

        $display("Test #1 Write 0xABCD to reg 0x5");
        axi_awaddr = 5'b00101 << 2;
        axi_wdata = 32'hABCD;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0011;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

        axi_arvalid = 1'b1;
        axi_araddr = 5'b00101 << 2;
        // Wait for AXI slave to send data
        wait (axi_arready == 1'b1);
        wait (axi_rvalid == 1'b1);
        assert (axi_rdata == 32'hABCD)
            $display("  - Read 0x%x value back successfully", axi_rdata);
        else
            $error("Failed to read correct value back, 0x%x != 0x%x", axi_rdata, 32'hABCD);
        // Signal to AXI Slave that data has been read
        axi_arvalid = 1'b0;
        axi_rready = 1'b1;
        wait (axi_rvalid == 1'b0);

        `reset_all
        $display("Test #1 Finished");

        $display("Test #2 Write 2 values, Read 2 values");
        $display("  - Writing 0xAAA0 to Reg 0");
        // Write to Reg #0
        axi_awaddr = 5'b00000 << 2;
        axi_wdata = 32'hAAA0;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0011;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

        // Write to Reg #1
        $display("  - Writing 0xAAA1 to Reg 1");
        axi_awaddr = 5'b00001 << 2;
        axi_wdata = 32'hAAA1;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0011;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

        $display("  - Now read both values back");
        // Read 1st value back
        axi_arvalid = 1'b1;
        axi_araddr = 5'b00000 << 2;
        // Wait for AXI slave to send data
        wait (axi_arready == 1'b1);
        wait (axi_rvalid == 1'b1);
        assert (axi_rdata == 32'hAAA0)
            $display("  - Read 0x%x value back successfully from Reg 0", axi_rdata);
        else
            $error("Failed to read correct value back, 0x%x != 0x%x", axi_rdata, 32'hAAA0);
        // Signal to AXI Slave that data has been read
        axi_arvalid = 1'b0;
        axi_rready = 1'b1;
        wait (axi_rvalid == 1'b0);
        // Delay between next operation
        `reset_all
        #20;

        // Read 2nd value back
        axi_arvalid = 1'b1;
        axi_araddr = 5'b00001 << 2;
        // Wait for AXI slave to send data
        wait (axi_arready == 1'b1);
        wait (axi_rvalid == 1'b1);
        assert (axi_rdata == 32'hAAA1)
            $display("  - Read 0x%x value back successfully from Reg 1", axi_rdata);
        else
            $error("Failed to read correct value back, 0x%x != 0x%x", axi_rdata, 32'hAAA1);
        // Signal to AXI Slave that data has been read
        axi_arvalid = 1'b0;
        axi_rready = 1'b1;
        wait (axi_rvalid == 1'b0);
        `reset_all
        #20;

        $display("Test #2 Finished");

        $display("Test #3 Prepare for I2C Write");
        // Write Address of Device to Reg #1
        $display("  - Writing Address of Device 0xFE to Reg 0");
        axi_awaddr = 5'b00000 << 2;
        axi_wdata = 32'h00005B;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0111;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

        // Write Address of Device to Reg #1
        $display("  - Writing Register Address 0x00 Reg 1");
        axi_awaddr = 5'b00001 << 2;
        axi_wdata = 32'h000000;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0111;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

        // Write Num of Bytes to Reg #2
        $display("  - Writing Register Address 0x00 Reg 2");
        axi_awaddr = 5'b00010 << 2;
        axi_wdata = 32'h0000FF;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0111;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

//        // Registers should now read:
//        // slv_reg0 <= 0x5B
//        // slv_reg1 <= 0x00
//        // slv_reg2 <= 0x01
        // Write 0 to Reg 7 (0x0) (I2C WRITE)
        $display("  - Writing Start (0x88) to Reg 7");
        axi_awaddr = 5'b00111 << 2;
        axi_wdata = 32'h88;
        axi_awvalid = 1'b1;
        axi_wstrb = 4'b0001;
        axi_wvalid = 1'b1;
        // Wait for AXI slave to ACK
        wait (axi_awready == 1'b1 &&
              axi_wready == 1'b1);
        wait (axi_awready == 1'b0 &&
              axi_wready == 1'b0);
        axi_awvalid = 0;
        axi_wvalid = 0;
        wait (axi_bvalid == 1'b1);
        // Ack
        axi_bready = 1'b1;
        wait (axi_bvalid == 1'b0);
        axi_bready = 1'b0;
        // Delay between next operation
        #10;
        `reset_all

        wait (busy == 0);
        wait (busy == 1'b0);

        wait (scl_io == 1);

        // Start condition
        wait (sda_io == 0);
        wait (scl_io == 0);
        #100;
        
        // Read 1st Byte (Slave address + direction)
        // 1011 011 [ 0 ]
        tmp_result = 8'b00000000;
        for (int i=0; i < 8; i++)
            begin
                tmp_result = (tmp_result << 1) | sda_io;
                #2500;
            end
        $display("Value read: %x", tmp_result);

        // ACK 1st byte (Slave address + direction)
        sda_drive = 1;
        sda_tx = 0;

        #2500;
        // Now slave releases the bus
        sda_drive = 0;

        // Read 2nd Byte (Register Address)
        // 0000 0000
        tmp_result = 8'b00000000;
        for (int i=0; i < 8; i++)
            begin
                tmp_result = (tmp_result << 1) | sda_io;
//                $display("bit #%d = %d", i, sda_io);
                #2500;
            end
        $display("Value read: %x", tmp_result);
        // ACK 2nd byte (Register Address)
        sda_drive = 1;
        sda_tx = 0;
        #2500;
        sda_drive = 0;

        // Read 3rd Byte (Value)
        tmp_result = 8'b00000000;
        for (int i=0; i < 8; i++)
            begin
                tmp_result = (tmp_result << 1) | sda_io;
//                $display("bit #%d = %d", i, sda_io);
                #2500;
            end
        $display("Value read: %x", tmp_result);
        // ACK 3rd byte (Value)
        sda_drive = 1;
        sda_tx = 0;
        #2500;
        sda_drive = 0;

        // STOP Condition
        wait (scl_io == 1);
        wait (sda_io == 1);
        // (Again?) Read 8 bits for Value

        #(2500 * 10);
        // Now initiate Read

        $display("  - Read Value from Reg 7");
        // Read Reg 7 (I2C READ)
        // Do a read on address 0x0
//        `reset_all
// JOHN
        axi_arvalid = 1'b1;
        axi_araddr = 5'b00111 << 2;
        // Wait for AXI slave to send data
        wait (axi_arready == 1'b1);
        wait (axi_rvalid == 1'b1);
        assert (axi_rdata == 32'hAAA1)
            $display("  - Read 0x%x value back successfully from Reg 1", axi_rdata);
        else
            $error("Failed to read correct value back, 0x%x != 0x%x", axi_rdata, 32'hAAA1);
        // Signal to AXI Slave that data has been read
        axi_arvalid = 1'b0;
        axi_rready = 1'b1;
        wait (axi_rvalid == 1'b0);
        `reset_all
        #20;

        $finish();




    end

    // Instantiate my_i2c_wrapper_v1_0_S00_AXI
    my_i2c_ip_v1_0_S00_AXI #(
        .C_S_AXI_DATA_WIDTH(32),
        .C_S_AXI_ADDR_WIDTH(5)
    )
        my_i2c_ip_dut(
            .scl_io(scl_io),
            .sda_io(sda_io),
            .req_data_chunk(req_data_chunk),
            .busy(busy),
            .nack(nack),
            // Global Clock Signal
            .S_AXI_ACLK(clk),

             //Global Reset Signal. This Signal is Active LOW
            .S_AXI_ARESETN(axi_aresetn),

            // Write address (issued by master, acceped by Slave)
            .S_AXI_AWADDR(axi_awaddr),

            // Write channel Protection type. This signal indicates the
    		// privilege and security level of the transaction, and whether
    		// the transaction is a data access or an instruction access.
            .S_AXI_AWPROT(axi_awprot),

            // Write address valid. This signal indicates that the master signaling
    		// valid write address and control information.
    		.S_AXI_AWVALID(axi_awvalid),

    		// Write address ready. This signal indicates that the slave is ready
    		// to accept an address and associated control signals.
            .S_AXI_AWREADY(axi_awready),

    		// Write data (issued by master, acceped by Slave) 
            .S_AXI_WDATA(axi_wdata),

            // Write strobes. This signal indicates which byte lanes hold
    		// valid data. There is one write strobe bit for each eight
    		// bits of the write data bus.    
            .S_AXI_WSTRB(axi_wstrb),

            // Write valid. This signal indicates that valid write
    		// data and strobes are available.
            .S_AXI_WVALID(axi_wvalid),

            // Write ready. This signal indicates that the slave
    		// can accept the write data.
		      .S_AXI_WREADY(axi_wready),

            // Write response. This signal indicates the status
    		// of the write transaction.
            .S_AXI_BRESP(axi_bresp),

    		// Write response valid. This signal indicates that the channel
    		// is signaling a valid write response.
            .S_AXI_BVALID(axi_bvalid),

            // Response ready. This signal indicates that the master
    		// can accept a write response.
		    .S_AXI_BREADY(axi_bready),

            // Read address (issued by master, acceped by Slave)
            .S_AXI_ARADDR(axi_araddr),

    		// Protection type. This signal indicates the privilege
    		// and security level of the transaction, and whether the
    		// transaction is a data access or an instruction access.
            .S_AXI_ARPROT(axi_arprot),

    		// Read address valid. This signal indicates that the channel
    		// is signaling valid read address and control information.
            .S_AXI_ARVALID(axi_arvalid),

            // Read address ready. This signal indicates that the slave is
    		// ready to accept an address and associated control signals.
            .S_AXI_ARREADY(axi_arready),

            // Read data (issued by slave)
            .S_AXI_RDATA(axi_rdata),

            // Read response. This signal indicates the status of the
    		// read transfer.
            .S_AXI_RRESP(axi_rresp),

            // Read valid. This signal indicates that the channel is
    		// signaling the required read data.
            .S_AXI_RVALID(axi_rvalid),

    		// Read ready. This signal indicates that the master can
    		// accept the read data and response information.
            .S_AXI_RREADY(axi_rready)
        );
endmodule
